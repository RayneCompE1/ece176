module helloVerilog ();

initial  
  $display("Hello Verilog!");

endmodule
