module s_decoder(input [3:0] i_bus, output reg [9:0] o_bus);

always @(*) 
begin
case (i_bus)
4'b0000: o_bus <= 10'b0000111111;
4'b0001: o_bus <= 10'b0000000110;
4'b0010: o_bus <= 10'b0001011011;
4'b0011: o_bus <= 10'b0001001111;
4'b0100: o_bus <= 10'b0001100110;
4'b0101: o_bus <= 10'b0001101101;
4'b0110: o_bus <= 10'b0001011111;
4'b0111: o_bus <= 10'b0000000111;
4'b1000: o_bus <= 10'b1001111111;
4'b1001: o_bus <= 10'b1000000111;
4'b1010: o_bus <= 10'b1001011111;
4'b1011: o_bus <= 10'b1001101101;
4'b1100: o_bus <= 10'b1001100110;
4'b1101: o_bus <= 10'b1001001111;
4'b1110: o_bus <= 10'b1001011011;
4'b1111: o_bus <= 10'b1000000110;
default: o_bus <= 10'b1111111111;
endcase
end

endmodule
